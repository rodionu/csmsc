-- MIPS Processor VHDL Behavioral Model
--
-- Ifetch module (provides the PC and instruction memory) 
-- 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Ifetch IS
	PORT(	SIGNAL Instruction 		: OUT	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
      		SIGNAL PC_OUT 			: OUT	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			SIGNAL PC_IN			: IN	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        	SIGNAL clock, reset 	: IN 	STD_LOGIC);
END Ifetch;

ARCHITECTURE behavior OF Ifetch IS
   TYPE INST_MEM IS ARRAY (0 to 18) of STD_LOGIC_VECTOR (31 DOWNTO 0);
   SIGNAL iram : INST_MEM := (
		X"3C011001",
		X"34280000",
		X"8D090000",
		X"8D0A0004",
		X"00001020",
		X"00006820",
		X"20030004",
		X"314C0001",
		X"34010000",
		X"102C0003",
		X"20630001",
		X"00491020",
		X"000A5042",
		X"00094840",
		X"21AD0001",
		X"20630008",
		X"34010010",
		X"142DFFF6",
		X"20630002"
   );
    
	SIGNAL PC	  			: STD_LOGIC_VECTOR( 31 DOWNTO 0 );
	SIGNAL Mem_Addr 		: STD_LOGIC_VECTOR( 31 DOWNTO 0 );
BEGIN 				
	--	PC(1 DOWNTO 0) <= "00";		
		PC_OUT <= PC;
  		Instruction <= iram(CONV_INTEGER(PC(31 DOWNTO 2)- X"0100000"));
	PROCESS
		BEGIN
			WAIT UNTIL ( clock'EVENT ) AND ( clock = '1' );
			IF reset = '1' THEN
				   PC( 31 DOWNTO 0) <= X"00400000"-4;
			ELSE 
				   PC( 31 DOWNTO 0 ) <= PC_IN( 31 DOWNTO 2) & "00";
			END IF;
			
	END PROCESS;
END behavior;


